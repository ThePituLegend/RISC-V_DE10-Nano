// UAB_RV_System.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module UAB_RV_System (
		input  wire        clk_clk,             //           clk.clk
		output wire [7:0]  leds_export,         //          leds.export
		output wire [14:0] memory_mem_a,        //        memory.mem_a
		output wire [2:0]  memory_mem_ba,       //              .mem_ba
		output wire        memory_mem_ck,       //              .mem_ck
		output wire        memory_mem_ck_n,     //              .mem_ck_n
		output wire        memory_mem_cke,      //              .mem_cke
		output wire        memory_mem_cs_n,     //              .mem_cs_n
		output wire        memory_mem_ras_n,    //              .mem_ras_n
		output wire        memory_mem_cas_n,    //              .mem_cas_n
		output wire        memory_mem_we_n,     //              .mem_we_n
		output wire        memory_mem_reset_n,  //              .mem_reset_n
		inout  wire [31:0] memory_mem_dq,       //              .mem_dq
		inout  wire [3:0]  memory_mem_dqs,      //              .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,    //              .mem_dqs_n
		output wire        memory_mem_odt,      //              .mem_odt
		output wire [3:0]  memory_mem_dm,       //              .mem_dm
		input  wire        memory_oct_rzqin,    //              .oct_rzqin
		input  wire        uabchip_reset_reset  // uabchip_reset.reset
	);

	wire          mem_pll_outclk0_clk;                                      // mem_pll:outclk_0 -> [ddr3:hps_f2h_sdram0_clock_clk, mm_interconnect_0:mem_pll_outclk0_clk, rst_controller_001:clk]
	wire          ddr3_h2f_reset_reset;                                     // ddr3:h2f_reset_reset_n -> [mem_pll:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire    [1:0] uabchip_0_axi4_mem_master_awburst;                        // UABChip_0:axi4_mem_0_bits_aw_bits_burst -> mm_interconnect_0:UABChip_0_axi4_mem_master_awburst
	wire    [7:0] uabchip_0_axi4_mem_master_arlen;                          // UABChip_0:axi4_mem_0_bits_ar_bits_len -> mm_interconnect_0:UABChip_0_axi4_mem_master_arlen
	wire    [3:0] uabchip_0_axi4_mem_master_arqos;                          // UABChip_0:axi4_mem_0_bits_ar_bits_qos -> mm_interconnect_0:UABChip_0_axi4_mem_master_arqos
	wire    [3:0] uabchip_0_axi4_mem_master_wstrb;                          // UABChip_0:axi4_mem_0_bits_w_bits_strb -> mm_interconnect_0:UABChip_0_axi4_mem_master_wstrb
	wire          uabchip_0_axi4_mem_master_wready;                         // mm_interconnect_0:UABChip_0_axi4_mem_master_wready -> UABChip_0:axi4_mem_0_bits_w_ready
	wire    [3:0] uabchip_0_axi4_mem_master_rid;                            // mm_interconnect_0:UABChip_0_axi4_mem_master_rid -> UABChip_0:axi4_mem_0_bits_r_bits_id
	wire          uabchip_0_axi4_mem_master_rready;                         // UABChip_0:axi4_mem_0_bits_r_ready -> mm_interconnect_0:UABChip_0_axi4_mem_master_rready
	wire    [7:0] uabchip_0_axi4_mem_master_awlen;                          // UABChip_0:axi4_mem_0_bits_aw_bits_len -> mm_interconnect_0:UABChip_0_axi4_mem_master_awlen
	wire    [3:0] uabchip_0_axi4_mem_master_awqos;                          // UABChip_0:axi4_mem_0_bits_aw_bits_qos -> mm_interconnect_0:UABChip_0_axi4_mem_master_awqos
	wire    [3:0] uabchip_0_axi4_mem_master_arcache;                        // UABChip_0:axi4_mem_0_bits_ar_bits_cache -> mm_interconnect_0:UABChip_0_axi4_mem_master_arcache
	wire   [31:0] uabchip_0_axi4_mem_master_araddr;                         // UABChip_0:axi4_mem_0_bits_ar_bits_addr -> mm_interconnect_0:UABChip_0_axi4_mem_master_araddr
	wire          uabchip_0_axi4_mem_master_wvalid;                         // UABChip_0:axi4_mem_0_bits_w_valid -> mm_interconnect_0:UABChip_0_axi4_mem_master_wvalid
	wire    [2:0] uabchip_0_axi4_mem_master_arprot;                         // UABChip_0:axi4_mem_0_bits_ar_bits_prot -> mm_interconnect_0:UABChip_0_axi4_mem_master_arprot
	wire          uabchip_0_axi4_mem_master_arvalid;                        // UABChip_0:axi4_mem_0_bits_ar_valid -> mm_interconnect_0:UABChip_0_axi4_mem_master_arvalid
	wire    [2:0] uabchip_0_axi4_mem_master_awprot;                         // UABChip_0:axi4_mem_0_bits_aw_bits_prot -> mm_interconnect_0:UABChip_0_axi4_mem_master_awprot
	wire   [31:0] uabchip_0_axi4_mem_master_wdata;                          // UABChip_0:axi4_mem_0_bits_w_bits_data -> mm_interconnect_0:UABChip_0_axi4_mem_master_wdata
	wire    [3:0] uabchip_0_axi4_mem_master_arid;                           // UABChip_0:axi4_mem_0_bits_ar_bits_id -> mm_interconnect_0:UABChip_0_axi4_mem_master_arid
	wire    [3:0] uabchip_0_axi4_mem_master_awcache;                        // UABChip_0:axi4_mem_0_bits_aw_bits_cache -> mm_interconnect_0:UABChip_0_axi4_mem_master_awcache
	wire          uabchip_0_axi4_mem_master_arlock;                         // UABChip_0:axi4_mem_0_bits_ar_bits_lock -> mm_interconnect_0:UABChip_0_axi4_mem_master_arlock
	wire          uabchip_0_axi4_mem_master_awlock;                         // UABChip_0:axi4_mem_0_bits_aw_bits_lock -> mm_interconnect_0:UABChip_0_axi4_mem_master_awlock
	wire   [31:0] uabchip_0_axi4_mem_master_awaddr;                         // UABChip_0:axi4_mem_0_bits_aw_bits_addr -> mm_interconnect_0:UABChip_0_axi4_mem_master_awaddr
	wire          uabchip_0_axi4_mem_master_arready;                        // mm_interconnect_0:UABChip_0_axi4_mem_master_arready -> UABChip_0:axi4_mem_0_bits_ar_ready
	wire    [1:0] uabchip_0_axi4_mem_master_bresp;                          // mm_interconnect_0:UABChip_0_axi4_mem_master_bresp -> UABChip_0:axi4_mem_0_bits_b_bits_resp
	wire   [31:0] uabchip_0_axi4_mem_master_rdata;                          // mm_interconnect_0:UABChip_0_axi4_mem_master_rdata -> UABChip_0:axi4_mem_0_bits_r_bits_data
	wire    [1:0] uabchip_0_axi4_mem_master_arburst;                        // UABChip_0:axi4_mem_0_bits_ar_bits_burst -> mm_interconnect_0:UABChip_0_axi4_mem_master_arburst
	wire          uabchip_0_axi4_mem_master_awready;                        // mm_interconnect_0:UABChip_0_axi4_mem_master_awready -> UABChip_0:axi4_mem_0_bits_aw_ready
	wire    [2:0] uabchip_0_axi4_mem_master_arsize;                         // UABChip_0:axi4_mem_0_bits_ar_bits_size -> mm_interconnect_0:UABChip_0_axi4_mem_master_arsize
	wire          uabchip_0_axi4_mem_master_bready;                         // UABChip_0:axi4_mem_0_bits_b_ready -> mm_interconnect_0:UABChip_0_axi4_mem_master_bready
	wire          uabchip_0_axi4_mem_master_rlast;                          // mm_interconnect_0:UABChip_0_axi4_mem_master_rlast -> UABChip_0:axi4_mem_0_bits_r_bits_last
	wire          uabchip_0_axi4_mem_master_wlast;                          // UABChip_0:axi4_mem_0_bits_w_bits_last -> mm_interconnect_0:UABChip_0_axi4_mem_master_wlast
	wire    [1:0] uabchip_0_axi4_mem_master_rresp;                          // mm_interconnect_0:UABChip_0_axi4_mem_master_rresp -> UABChip_0:axi4_mem_0_bits_r_bits_resp
	wire    [3:0] uabchip_0_axi4_mem_master_awid;                           // UABChip_0:axi4_mem_0_bits_aw_bits_id -> mm_interconnect_0:UABChip_0_axi4_mem_master_awid
	wire    [3:0] uabchip_0_axi4_mem_master_bid;                            // mm_interconnect_0:UABChip_0_axi4_mem_master_bid -> UABChip_0:axi4_mem_0_bits_b_bits_id
	wire          uabchip_0_axi4_mem_master_bvalid;                         // mm_interconnect_0:UABChip_0_axi4_mem_master_bvalid -> UABChip_0:axi4_mem_0_bits_b_valid
	wire    [2:0] uabchip_0_axi4_mem_master_awsize;                         // UABChip_0:axi4_mem_0_bits_aw_bits_size -> mm_interconnect_0:UABChip_0_axi4_mem_master_awsize
	wire          uabchip_0_axi4_mem_master_awvalid;                        // UABChip_0:axi4_mem_0_bits_aw_valid -> mm_interconnect_0:UABChip_0_axi4_mem_master_awvalid
	wire          uabchip_0_axi4_mem_master_rvalid;                         // mm_interconnect_0:UABChip_0_axi4_mem_master_rvalid -> UABChip_0:axi4_mem_0_bits_r_valid
	wire  [127:0] mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdata;      // ddr3:hps_f2h_sdram0_data_readdata -> mm_interconnect_0:ddr3_hps_f2h_sdram0_data_readdata
	wire          mm_interconnect_0_ddr3_hps_f2h_sdram0_data_waitrequest;   // ddr3:hps_f2h_sdram0_data_waitrequest -> mm_interconnect_0:ddr3_hps_f2h_sdram0_data_waitrequest
	wire   [25:0] mm_interconnect_0_ddr3_hps_f2h_sdram0_data_address;       // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_address -> ddr3:hps_f2h_sdram0_data_address
	wire          mm_interconnect_0_ddr3_hps_f2h_sdram0_data_read;          // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_read -> ddr3:hps_f2h_sdram0_data_read
	wire   [15:0] mm_interconnect_0_ddr3_hps_f2h_sdram0_data_byteenable;    // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_byteenable -> ddr3:hps_f2h_sdram0_data_byteenable
	wire          mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdatavalid; // ddr3:hps_f2h_sdram0_data_readdatavalid -> mm_interconnect_0:ddr3_hps_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_0_ddr3_hps_f2h_sdram0_data_write;         // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_write -> ddr3:hps_f2h_sdram0_data_write
	wire  [127:0] mm_interconnect_0_ddr3_hps_f2h_sdram0_data_writedata;     // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_writedata -> ddr3:hps_f2h_sdram0_data_writedata
	wire    [8:0] mm_interconnect_0_ddr3_hps_f2h_sdram0_data_burstcount;    // mm_interconnect_0:ddr3_hps_f2h_sdram0_data_burstcount -> ddr3:hps_f2h_sdram0_data_burstcount
	wire    [1:0] uabchip_0_axi4_mmio_master_awburst;                       // UABChip_0:axi4_mmio_0_bits_aw_bits_burst -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awburst
	wire    [7:0] uabchip_0_axi4_mmio_master_arlen;                         // UABChip_0:axi4_mmio_0_bits_ar_bits_len -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arlen
	wire    [3:0] uabchip_0_axi4_mmio_master_arqos;                         // UABChip_0:axi4_mmio_0_bits_ar_bits_qos -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arqos
	wire    [3:0] uabchip_0_axi4_mmio_master_wstrb;                         // UABChip_0:axi4_mmio_0_bits_w_bits_strb -> mm_interconnect_1:UABChip_0_axi4_mmio_master_wstrb
	wire          uabchip_0_axi4_mmio_master_wready;                        // mm_interconnect_1:UABChip_0_axi4_mmio_master_wready -> UABChip_0:axi4_mmio_0_bits_w_ready
	wire    [3:0] uabchip_0_axi4_mmio_master_rid;                           // mm_interconnect_1:UABChip_0_axi4_mmio_master_rid -> UABChip_0:axi4_mmio_0_bits_r_bits_id
	wire          uabchip_0_axi4_mmio_master_rready;                        // UABChip_0:axi4_mmio_0_bits_r_ready -> mm_interconnect_1:UABChip_0_axi4_mmio_master_rready
	wire    [7:0] uabchip_0_axi4_mmio_master_awlen;                         // UABChip_0:axi4_mmio_0_bits_aw_bits_len -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awlen
	wire    [3:0] uabchip_0_axi4_mmio_master_awqos;                         // UABChip_0:axi4_mmio_0_bits_aw_bits_qos -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awqos
	wire    [3:0] uabchip_0_axi4_mmio_master_arcache;                       // UABChip_0:axi4_mmio_0_bits_ar_bits_cache -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arcache
	wire   [30:0] uabchip_0_axi4_mmio_master_araddr;                        // UABChip_0:axi4_mmio_0_bits_ar_bits_addr -> mm_interconnect_1:UABChip_0_axi4_mmio_master_araddr
	wire          uabchip_0_axi4_mmio_master_wvalid;                        // UABChip_0:axi4_mmio_0_bits_w_valid -> mm_interconnect_1:UABChip_0_axi4_mmio_master_wvalid
	wire    [2:0] uabchip_0_axi4_mmio_master_arprot;                        // UABChip_0:axi4_mmio_0_bits_ar_bits_prot -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arprot
	wire          uabchip_0_axi4_mmio_master_arvalid;                       // UABChip_0:axi4_mmio_0_bits_ar_valid -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arvalid
	wire    [2:0] uabchip_0_axi4_mmio_master_awprot;                        // UABChip_0:axi4_mmio_0_bits_aw_bits_prot -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awprot
	wire   [31:0] uabchip_0_axi4_mmio_master_wdata;                         // UABChip_0:axi4_mmio_0_bits_w_bits_data -> mm_interconnect_1:UABChip_0_axi4_mmio_master_wdata
	wire    [3:0] uabchip_0_axi4_mmio_master_arid;                          // UABChip_0:axi4_mmio_0_bits_ar_bits_id -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arid
	wire    [3:0] uabchip_0_axi4_mmio_master_awcache;                       // UABChip_0:axi4_mmio_0_bits_aw_bits_cache -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awcache
	wire          uabchip_0_axi4_mmio_master_arlock;                        // UABChip_0:axi4_mmio_0_bits_ar_bits_lock -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arlock
	wire          uabchip_0_axi4_mmio_master_awlock;                        // UABChip_0:axi4_mmio_0_bits_aw_bits_lock -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awlock
	wire   [30:0] uabchip_0_axi4_mmio_master_awaddr;                        // UABChip_0:axi4_mmio_0_bits_aw_bits_addr -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awaddr
	wire          uabchip_0_axi4_mmio_master_arready;                       // mm_interconnect_1:UABChip_0_axi4_mmio_master_arready -> UABChip_0:axi4_mmio_0_bits_ar_ready
	wire    [1:0] uabchip_0_axi4_mmio_master_bresp;                         // mm_interconnect_1:UABChip_0_axi4_mmio_master_bresp -> UABChip_0:axi4_mmio_0_bits_b_bits_resp
	wire   [31:0] uabchip_0_axi4_mmio_master_rdata;                         // mm_interconnect_1:UABChip_0_axi4_mmio_master_rdata -> UABChip_0:axi4_mmio_0_bits_r_bits_data
	wire    [1:0] uabchip_0_axi4_mmio_master_arburst;                       // UABChip_0:axi4_mmio_0_bits_ar_bits_burst -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arburst
	wire          uabchip_0_axi4_mmio_master_awready;                       // mm_interconnect_1:UABChip_0_axi4_mmio_master_awready -> UABChip_0:axi4_mmio_0_bits_aw_ready
	wire    [2:0] uabchip_0_axi4_mmio_master_arsize;                        // UABChip_0:axi4_mmio_0_bits_ar_bits_size -> mm_interconnect_1:UABChip_0_axi4_mmio_master_arsize
	wire          uabchip_0_axi4_mmio_master_bready;                        // UABChip_0:axi4_mmio_0_bits_b_ready -> mm_interconnect_1:UABChip_0_axi4_mmio_master_bready
	wire          uabchip_0_axi4_mmio_master_rlast;                         // mm_interconnect_1:UABChip_0_axi4_mmio_master_rlast -> UABChip_0:axi4_mmio_0_bits_r_bits_last
	wire          uabchip_0_axi4_mmio_master_wlast;                         // UABChip_0:axi4_mmio_0_bits_w_bits_last -> mm_interconnect_1:UABChip_0_axi4_mmio_master_wlast
	wire    [1:0] uabchip_0_axi4_mmio_master_rresp;                         // mm_interconnect_1:UABChip_0_axi4_mmio_master_rresp -> UABChip_0:axi4_mmio_0_bits_r_bits_resp
	wire    [3:0] uabchip_0_axi4_mmio_master_awid;                          // UABChip_0:axi4_mmio_0_bits_aw_bits_id -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awid
	wire    [3:0] uabchip_0_axi4_mmio_master_bid;                           // mm_interconnect_1:UABChip_0_axi4_mmio_master_bid -> UABChip_0:axi4_mmio_0_bits_b_bits_id
	wire          uabchip_0_axi4_mmio_master_bvalid;                        // mm_interconnect_1:UABChip_0_axi4_mmio_master_bvalid -> UABChip_0:axi4_mmio_0_bits_b_valid
	wire    [2:0] uabchip_0_axi4_mmio_master_awsize;                        // UABChip_0:axi4_mmio_0_bits_aw_bits_size -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awsize
	wire          uabchip_0_axi4_mmio_master_awvalid;                       // UABChip_0:axi4_mmio_0_bits_aw_valid -> mm_interconnect_1:UABChip_0_axi4_mmio_master_awvalid
	wire          uabchip_0_axi4_mmio_master_rvalid;                        // mm_interconnect_1:UABChip_0_axi4_mmio_master_rvalid -> UABChip_0:axi4_mmio_0_bits_r_valid
	wire          mm_interconnect_1_onchip_memory_s1_chipselect;            // mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire   [63:0] mm_interconnect_1_onchip_memory_s1_readdata;              // onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	wire   [12:0] mm_interconnect_1_onchip_memory_s1_address;               // mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	wire    [7:0] mm_interconnect_1_onchip_memory_s1_byteenable;            // mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire          mm_interconnect_1_onchip_memory_s1_write;                 // mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	wire   [63:0] mm_interconnect_1_onchip_memory_s1_writedata;             // mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire          mm_interconnect_1_onchip_memory_s1_clken;                 // mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	wire          mm_interconnect_1_pio_0_s1_chipselect;                    // mm_interconnect_1:pio_0_s1_chipselect -> pio_0:chipselect
	wire   [31:0] mm_interconnect_1_pio_0_s1_readdata;                      // pio_0:readdata -> mm_interconnect_1:pio_0_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_0_s1_address;                       // mm_interconnect_1:pio_0_s1_address -> pio_0:address
	wire          mm_interconnect_1_pio_0_s1_write;                         // mm_interconnect_1:pio_0_s1_write -> pio_0:write_n
	wire   [31:0] mm_interconnect_1_pio_0_s1_writedata;                     // mm_interconnect_1:pio_0_s1_writedata -> pio_0:writedata
	wire          rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [mm_interconnect_1:onchip_memory_reset1_reset_bridge_in_reset_reset, onchip_memory:reset, pio_0:reset_n]
	wire          rst_controller_reset_out_reset_req;                       // rst_controller:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> mm_interconnect_0:ddr3_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset

	ChipTop uabchip_0 (
		.clock                          (clk_clk),                            //            clock.clk
		.reset_wire_reset               (uabchip_reset_reset),                //            reset.reset
		.axi4_mem_0_bits_ar_bits_addr   (uabchip_0_axi4_mem_master_araddr),   //  axi4_mem_master.araddr
		.axi4_mem_0_bits_ar_bits_burst  (uabchip_0_axi4_mem_master_arburst),  //                 .arburst
		.axi4_mem_0_bits_ar_bits_cache  (uabchip_0_axi4_mem_master_arcache),  //                 .arcache
		.axi4_mem_0_bits_ar_bits_id     (uabchip_0_axi4_mem_master_arid),     //                 .arid
		.axi4_mem_0_bits_ar_bits_len    (uabchip_0_axi4_mem_master_arlen),    //                 .arlen
		.axi4_mem_0_bits_ar_bits_lock   (uabchip_0_axi4_mem_master_arlock),   //                 .arlock
		.axi4_mem_0_bits_ar_bits_prot   (uabchip_0_axi4_mem_master_arprot),   //                 .arprot
		.axi4_mem_0_bits_ar_bits_qos    (uabchip_0_axi4_mem_master_arqos),    //                 .arqos
		.axi4_mem_0_bits_ar_bits_size   (uabchip_0_axi4_mem_master_arsize),   //                 .arsize
		.axi4_mem_0_bits_ar_ready       (uabchip_0_axi4_mem_master_arready),  //                 .arready
		.axi4_mem_0_bits_ar_valid       (uabchip_0_axi4_mem_master_arvalid),  //                 .arvalid
		.axi4_mem_0_bits_aw_bits_addr   (uabchip_0_axi4_mem_master_awaddr),   //                 .awaddr
		.axi4_mem_0_bits_aw_bits_burst  (uabchip_0_axi4_mem_master_awburst),  //                 .awburst
		.axi4_mem_0_bits_aw_bits_cache  (uabchip_0_axi4_mem_master_awcache),  //                 .awcache
		.axi4_mem_0_bits_aw_bits_id     (uabchip_0_axi4_mem_master_awid),     //                 .awid
		.axi4_mem_0_bits_aw_bits_len    (uabchip_0_axi4_mem_master_awlen),    //                 .awlen
		.axi4_mem_0_bits_aw_bits_lock   (uabchip_0_axi4_mem_master_awlock),   //                 .awlock
		.axi4_mem_0_bits_aw_bits_prot   (uabchip_0_axi4_mem_master_awprot),   //                 .awprot
		.axi4_mem_0_bits_aw_bits_qos    (uabchip_0_axi4_mem_master_awqos),    //                 .awqos
		.axi4_mem_0_bits_aw_bits_size   (uabchip_0_axi4_mem_master_awsize),   //                 .awsize
		.axi4_mem_0_bits_aw_ready       (uabchip_0_axi4_mem_master_awready),  //                 .awready
		.axi4_mem_0_bits_aw_valid       (uabchip_0_axi4_mem_master_awvalid),  //                 .awvalid
		.axi4_mem_0_bits_b_bits_id      (uabchip_0_axi4_mem_master_bid),      //                 .bid
		.axi4_mem_0_bits_b_bits_resp    (uabchip_0_axi4_mem_master_bresp),    //                 .bresp
		.axi4_mem_0_bits_b_ready        (uabchip_0_axi4_mem_master_bready),   //                 .bready
		.axi4_mem_0_bits_b_valid        (uabchip_0_axi4_mem_master_bvalid),   //                 .bvalid
		.axi4_mem_0_bits_r_bits_data    (uabchip_0_axi4_mem_master_rdata),    //                 .rdata
		.axi4_mem_0_bits_r_bits_id      (uabchip_0_axi4_mem_master_rid),      //                 .rid
		.axi4_mem_0_bits_r_bits_last    (uabchip_0_axi4_mem_master_rlast),    //                 .rlast
		.axi4_mem_0_bits_r_bits_resp    (uabchip_0_axi4_mem_master_rresp),    //                 .rresp
		.axi4_mem_0_bits_r_ready        (uabchip_0_axi4_mem_master_rready),   //                 .rready
		.axi4_mem_0_bits_r_valid        (uabchip_0_axi4_mem_master_rvalid),   //                 .rvalid
		.axi4_mem_0_bits_w_bits_data    (uabchip_0_axi4_mem_master_wdata),    //                 .wdata
		.axi4_mem_0_bits_w_bits_last    (uabchip_0_axi4_mem_master_wlast),    //                 .wlast
		.axi4_mem_0_bits_w_bits_strb    (uabchip_0_axi4_mem_master_wstrb),    //                 .wstrb
		.axi4_mem_0_bits_w_ready        (uabchip_0_axi4_mem_master_wready),   //                 .wready
		.axi4_mem_0_bits_w_valid        (uabchip_0_axi4_mem_master_wvalid),   //                 .wvalid
		.axi4_mmio_0_bits_ar_bits_addr  (uabchip_0_axi4_mmio_master_araddr),  // axi4_mmio_master.araddr
		.axi4_mmio_0_bits_ar_bits_burst (uabchip_0_axi4_mmio_master_arburst), //                 .arburst
		.axi4_mmio_0_bits_ar_bits_cache (uabchip_0_axi4_mmio_master_arcache), //                 .arcache
		.axi4_mmio_0_bits_ar_bits_id    (uabchip_0_axi4_mmio_master_arid),    //                 .arid
		.axi4_mmio_0_bits_ar_bits_len   (uabchip_0_axi4_mmio_master_arlen),   //                 .arlen
		.axi4_mmio_0_bits_ar_bits_lock  (uabchip_0_axi4_mmio_master_arlock),  //                 .arlock
		.axi4_mmio_0_bits_ar_bits_prot  (uabchip_0_axi4_mmio_master_arprot),  //                 .arprot
		.axi4_mmio_0_bits_ar_bits_qos   (uabchip_0_axi4_mmio_master_arqos),   //                 .arqos
		.axi4_mmio_0_bits_ar_bits_size  (uabchip_0_axi4_mmio_master_arsize),  //                 .arsize
		.axi4_mmio_0_bits_ar_ready      (uabchip_0_axi4_mmio_master_arready), //                 .arready
		.axi4_mmio_0_bits_ar_valid      (uabchip_0_axi4_mmio_master_arvalid), //                 .arvalid
		.axi4_mmio_0_bits_aw_bits_addr  (uabchip_0_axi4_mmio_master_awaddr),  //                 .awaddr
		.axi4_mmio_0_bits_aw_bits_burst (uabchip_0_axi4_mmio_master_awburst), //                 .awburst
		.axi4_mmio_0_bits_aw_bits_cache (uabchip_0_axi4_mmio_master_awcache), //                 .awcache
		.axi4_mmio_0_bits_aw_bits_id    (uabchip_0_axi4_mmio_master_awid),    //                 .awid
		.axi4_mmio_0_bits_aw_bits_len   (uabchip_0_axi4_mmio_master_awlen),   //                 .awlen
		.axi4_mmio_0_bits_aw_bits_lock  (uabchip_0_axi4_mmio_master_awlock),  //                 .awlock
		.axi4_mmio_0_bits_aw_bits_prot  (uabchip_0_axi4_mmio_master_awprot),  //                 .awprot
		.axi4_mmio_0_bits_aw_bits_qos   (uabchip_0_axi4_mmio_master_awqos),   //                 .awqos
		.axi4_mmio_0_bits_aw_bits_size  (uabchip_0_axi4_mmio_master_awsize),  //                 .awsize
		.axi4_mmio_0_bits_aw_ready      (uabchip_0_axi4_mmio_master_awready), //                 .awready
		.axi4_mmio_0_bits_aw_valid      (uabchip_0_axi4_mmio_master_awvalid), //                 .awvalid
		.axi4_mmio_0_bits_b_bits_id     (uabchip_0_axi4_mmio_master_bid),     //                 .bid
		.axi4_mmio_0_bits_b_bits_resp   (uabchip_0_axi4_mmio_master_bresp),   //                 .bresp
		.axi4_mmio_0_bits_b_ready       (uabchip_0_axi4_mmio_master_bready),  //                 .bready
		.axi4_mmio_0_bits_b_valid       (uabchip_0_axi4_mmio_master_bvalid),  //                 .bvalid
		.axi4_mmio_0_bits_r_bits_data   (uabchip_0_axi4_mmio_master_rdata),   //                 .rdata
		.axi4_mmio_0_bits_r_bits_id     (uabchip_0_axi4_mmio_master_rid),     //                 .rid
		.axi4_mmio_0_bits_r_bits_last   (uabchip_0_axi4_mmio_master_rlast),   //                 .rlast
		.axi4_mmio_0_bits_r_bits_resp   (uabchip_0_axi4_mmio_master_rresp),   //                 .rresp
		.axi4_mmio_0_bits_r_ready       (uabchip_0_axi4_mmio_master_rready),  //                 .rready
		.axi4_mmio_0_bits_r_valid       (uabchip_0_axi4_mmio_master_rvalid),  //                 .rvalid
		.axi4_mmio_0_bits_w_bits_data   (uabchip_0_axi4_mmio_master_wdata),   //                 .wdata
		.axi4_mmio_0_bits_w_bits_last   (uabchip_0_axi4_mmio_master_wlast),   //                 .wlast
		.axi4_mmio_0_bits_w_bits_strb   (uabchip_0_axi4_mmio_master_wstrb),   //                 .wstrb
		.axi4_mmio_0_bits_w_ready       (uabchip_0_axi4_mmio_master_wready),  //                 .wready
		.axi4_mmio_0_bits_w_valid       (uabchip_0_axi4_mmio_master_wvalid)   //                 .wvalid
	);

	UAB_RV_System_ddr3 ddr3 (
		.clk_clk                           (clk_clk),                                                  //                  clk.clk
		.h2f_reset_reset_n                 (ddr3_h2f_reset_reset),                                     //            h2f_reset.reset_n
		.hps_f2h_sdram0_clock_clk          (mem_pll_outclk0_clk),                                      // hps_f2h_sdram0_clock.clk
		.hps_f2h_sdram0_data_address       (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_address),       //  hps_f2h_sdram0_data.address
		.hps_f2h_sdram0_data_read          (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_read),          //                     .read
		.hps_f2h_sdram0_data_readdata      (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdata),      //                     .readdata
		.hps_f2h_sdram0_data_write         (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_write),         //                     .write
		.hps_f2h_sdram0_data_writedata     (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_writedata),     //                     .writedata
		.hps_f2h_sdram0_data_readdatavalid (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdatavalid), //                     .readdatavalid
		.hps_f2h_sdram0_data_waitrequest   (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_waitrequest),   //                     .waitrequest
		.hps_f2h_sdram0_data_byteenable    (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_byteenable),    //                     .byteenable
		.hps_f2h_sdram0_data_burstcount    (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_burstcount),    //                     .burstcount
		.memory_mem_a                      (memory_mem_a),                                             //               memory.mem_a
		.memory_mem_ba                     (memory_mem_ba),                                            //                     .mem_ba
		.memory_mem_ck                     (memory_mem_ck),                                            //                     .mem_ck
		.memory_mem_ck_n                   (memory_mem_ck_n),                                          //                     .mem_ck_n
		.memory_mem_cke                    (memory_mem_cke),                                           //                     .mem_cke
		.memory_mem_cs_n                   (memory_mem_cs_n),                                          //                     .mem_cs_n
		.memory_mem_ras_n                  (memory_mem_ras_n),                                         //                     .mem_ras_n
		.memory_mem_cas_n                  (memory_mem_cas_n),                                         //                     .mem_cas_n
		.memory_mem_we_n                   (memory_mem_we_n),                                          //                     .mem_we_n
		.memory_mem_reset_n                (memory_mem_reset_n),                                       //                     .mem_reset_n
		.memory_mem_dq                     (memory_mem_dq),                                            //                     .mem_dq
		.memory_mem_dqs                    (memory_mem_dqs),                                           //                     .mem_dqs
		.memory_mem_dqs_n                  (memory_mem_dqs_n),                                         //                     .mem_dqs_n
		.memory_mem_odt                    (memory_mem_odt),                                           //                     .mem_odt
		.memory_mem_dm                     (memory_mem_dm),                                            //                     .mem_dm
		.memory_oct_rzqin                  (memory_oct_rzqin)                                          //                     .oct_rzqin
	);

	UAB_RV_System_mem_pll mem_pll (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~ddr3_h2f_reset_reset), //   reset.reset
		.outclk_0 (mem_pll_outclk0_clk),   // outclk0.clk
		.locked   ()                       // (terminated)
	);

	UAB_RV_System_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	UAB_RV_System_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_1_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_0_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                            // external_connection.export
	);

	UAB_RV_System_mm_interconnect_0 mm_interconnect_0 (
		.UABChip_0_axi4_mem_master_awid                                        (uabchip_0_axi4_mem_master_awid),                           //                                       UABChip_0_axi4_mem_master.awid
		.UABChip_0_axi4_mem_master_awaddr                                      (uabchip_0_axi4_mem_master_awaddr),                         //                                                                .awaddr
		.UABChip_0_axi4_mem_master_awlen                                       (uabchip_0_axi4_mem_master_awlen),                          //                                                                .awlen
		.UABChip_0_axi4_mem_master_awsize                                      (uabchip_0_axi4_mem_master_awsize),                         //                                                                .awsize
		.UABChip_0_axi4_mem_master_awburst                                     (uabchip_0_axi4_mem_master_awburst),                        //                                                                .awburst
		.UABChip_0_axi4_mem_master_awlock                                      (uabchip_0_axi4_mem_master_awlock),                         //                                                                .awlock
		.UABChip_0_axi4_mem_master_awcache                                     (uabchip_0_axi4_mem_master_awcache),                        //                                                                .awcache
		.UABChip_0_axi4_mem_master_awprot                                      (uabchip_0_axi4_mem_master_awprot),                         //                                                                .awprot
		.UABChip_0_axi4_mem_master_awqos                                       (uabchip_0_axi4_mem_master_awqos),                          //                                                                .awqos
		.UABChip_0_axi4_mem_master_awvalid                                     (uabchip_0_axi4_mem_master_awvalid),                        //                                                                .awvalid
		.UABChip_0_axi4_mem_master_awready                                     (uabchip_0_axi4_mem_master_awready),                        //                                                                .awready
		.UABChip_0_axi4_mem_master_wdata                                       (uabchip_0_axi4_mem_master_wdata),                          //                                                                .wdata
		.UABChip_0_axi4_mem_master_wstrb                                       (uabchip_0_axi4_mem_master_wstrb),                          //                                                                .wstrb
		.UABChip_0_axi4_mem_master_wlast                                       (uabchip_0_axi4_mem_master_wlast),                          //                                                                .wlast
		.UABChip_0_axi4_mem_master_wvalid                                      (uabchip_0_axi4_mem_master_wvalid),                         //                                                                .wvalid
		.UABChip_0_axi4_mem_master_wready                                      (uabchip_0_axi4_mem_master_wready),                         //                                                                .wready
		.UABChip_0_axi4_mem_master_bid                                         (uabchip_0_axi4_mem_master_bid),                            //                                                                .bid
		.UABChip_0_axi4_mem_master_bresp                                       (uabchip_0_axi4_mem_master_bresp),                          //                                                                .bresp
		.UABChip_0_axi4_mem_master_bvalid                                      (uabchip_0_axi4_mem_master_bvalid),                         //                                                                .bvalid
		.UABChip_0_axi4_mem_master_bready                                      (uabchip_0_axi4_mem_master_bready),                         //                                                                .bready
		.UABChip_0_axi4_mem_master_arid                                        (uabchip_0_axi4_mem_master_arid),                           //                                                                .arid
		.UABChip_0_axi4_mem_master_araddr                                      (uabchip_0_axi4_mem_master_araddr),                         //                                                                .araddr
		.UABChip_0_axi4_mem_master_arlen                                       (uabchip_0_axi4_mem_master_arlen),                          //                                                                .arlen
		.UABChip_0_axi4_mem_master_arsize                                      (uabchip_0_axi4_mem_master_arsize),                         //                                                                .arsize
		.UABChip_0_axi4_mem_master_arburst                                     (uabchip_0_axi4_mem_master_arburst),                        //                                                                .arburst
		.UABChip_0_axi4_mem_master_arlock                                      (uabchip_0_axi4_mem_master_arlock),                         //                                                                .arlock
		.UABChip_0_axi4_mem_master_arcache                                     (uabchip_0_axi4_mem_master_arcache),                        //                                                                .arcache
		.UABChip_0_axi4_mem_master_arprot                                      (uabchip_0_axi4_mem_master_arprot),                         //                                                                .arprot
		.UABChip_0_axi4_mem_master_arqos                                       (uabchip_0_axi4_mem_master_arqos),                          //                                                                .arqos
		.UABChip_0_axi4_mem_master_arvalid                                     (uabchip_0_axi4_mem_master_arvalid),                        //                                                                .arvalid
		.UABChip_0_axi4_mem_master_arready                                     (uabchip_0_axi4_mem_master_arready),                        //                                                                .arready
		.UABChip_0_axi4_mem_master_rid                                         (uabchip_0_axi4_mem_master_rid),                            //                                                                .rid
		.UABChip_0_axi4_mem_master_rdata                                       (uabchip_0_axi4_mem_master_rdata),                          //                                                                .rdata
		.UABChip_0_axi4_mem_master_rresp                                       (uabchip_0_axi4_mem_master_rresp),                          //                                                                .rresp
		.UABChip_0_axi4_mem_master_rlast                                       (uabchip_0_axi4_mem_master_rlast),                          //                                                                .rlast
		.UABChip_0_axi4_mem_master_rvalid                                      (uabchip_0_axi4_mem_master_rvalid),                         //                                                                .rvalid
		.UABChip_0_axi4_mem_master_rready                                      (uabchip_0_axi4_mem_master_rready),                         //                                                                .rready
		.clk_clk_clk                                                           (clk_clk),                                                  //                                                         clk_clk.clk
		.mem_pll_outclk0_clk                                                   (mem_pll_outclk0_clk),                                      //                                                 mem_pll_outclk0.clk
		.ddr3_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // ddr3_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.UABChip_0_reset_reset_bridge_in_reset_reset                           (uabchip_reset_reset),                                      //                           UABChip_0_reset_reset_bridge_in_reset.reset
		.ddr3_hps_f2h_sdram0_data_address                                      (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_address),       //                                        ddr3_hps_f2h_sdram0_data.address
		.ddr3_hps_f2h_sdram0_data_write                                        (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_write),         //                                                                .write
		.ddr3_hps_f2h_sdram0_data_read                                         (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_read),          //                                                                .read
		.ddr3_hps_f2h_sdram0_data_readdata                                     (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdata),      //                                                                .readdata
		.ddr3_hps_f2h_sdram0_data_writedata                                    (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_writedata),     //                                                                .writedata
		.ddr3_hps_f2h_sdram0_data_burstcount                                   (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_burstcount),    //                                                                .burstcount
		.ddr3_hps_f2h_sdram0_data_byteenable                                   (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_byteenable),    //                                                                .byteenable
		.ddr3_hps_f2h_sdram0_data_readdatavalid                                (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_readdatavalid), //                                                                .readdatavalid
		.ddr3_hps_f2h_sdram0_data_waitrequest                                  (mm_interconnect_0_ddr3_hps_f2h_sdram0_data_waitrequest)    //                                                                .waitrequest
	);

	UAB_RV_System_mm_interconnect_1 mm_interconnect_1 (
		.UABChip_0_axi4_mmio_master_awid                  (uabchip_0_axi4_mmio_master_awid),               //                 UABChip_0_axi4_mmio_master.awid
		.UABChip_0_axi4_mmio_master_awaddr                (uabchip_0_axi4_mmio_master_awaddr),             //                                           .awaddr
		.UABChip_0_axi4_mmio_master_awlen                 (uabchip_0_axi4_mmio_master_awlen),              //                                           .awlen
		.UABChip_0_axi4_mmio_master_awsize                (uabchip_0_axi4_mmio_master_awsize),             //                                           .awsize
		.UABChip_0_axi4_mmio_master_awburst               (uabchip_0_axi4_mmio_master_awburst),            //                                           .awburst
		.UABChip_0_axi4_mmio_master_awlock                (uabchip_0_axi4_mmio_master_awlock),             //                                           .awlock
		.UABChip_0_axi4_mmio_master_awcache               (uabchip_0_axi4_mmio_master_awcache),            //                                           .awcache
		.UABChip_0_axi4_mmio_master_awprot                (uabchip_0_axi4_mmio_master_awprot),             //                                           .awprot
		.UABChip_0_axi4_mmio_master_awqos                 (uabchip_0_axi4_mmio_master_awqos),              //                                           .awqos
		.UABChip_0_axi4_mmio_master_awvalid               (uabchip_0_axi4_mmio_master_awvalid),            //                                           .awvalid
		.UABChip_0_axi4_mmio_master_awready               (uabchip_0_axi4_mmio_master_awready),            //                                           .awready
		.UABChip_0_axi4_mmio_master_wdata                 (uabchip_0_axi4_mmio_master_wdata),              //                                           .wdata
		.UABChip_0_axi4_mmio_master_wstrb                 (uabchip_0_axi4_mmio_master_wstrb),              //                                           .wstrb
		.UABChip_0_axi4_mmio_master_wlast                 (uabchip_0_axi4_mmio_master_wlast),              //                                           .wlast
		.UABChip_0_axi4_mmio_master_wvalid                (uabchip_0_axi4_mmio_master_wvalid),             //                                           .wvalid
		.UABChip_0_axi4_mmio_master_wready                (uabchip_0_axi4_mmio_master_wready),             //                                           .wready
		.UABChip_0_axi4_mmio_master_bid                   (uabchip_0_axi4_mmio_master_bid),                //                                           .bid
		.UABChip_0_axi4_mmio_master_bresp                 (uabchip_0_axi4_mmio_master_bresp),              //                                           .bresp
		.UABChip_0_axi4_mmio_master_bvalid                (uabchip_0_axi4_mmio_master_bvalid),             //                                           .bvalid
		.UABChip_0_axi4_mmio_master_bready                (uabchip_0_axi4_mmio_master_bready),             //                                           .bready
		.UABChip_0_axi4_mmio_master_arid                  (uabchip_0_axi4_mmio_master_arid),               //                                           .arid
		.UABChip_0_axi4_mmio_master_araddr                (uabchip_0_axi4_mmio_master_araddr),             //                                           .araddr
		.UABChip_0_axi4_mmio_master_arlen                 (uabchip_0_axi4_mmio_master_arlen),              //                                           .arlen
		.UABChip_0_axi4_mmio_master_arsize                (uabchip_0_axi4_mmio_master_arsize),             //                                           .arsize
		.UABChip_0_axi4_mmio_master_arburst               (uabchip_0_axi4_mmio_master_arburst),            //                                           .arburst
		.UABChip_0_axi4_mmio_master_arlock                (uabchip_0_axi4_mmio_master_arlock),             //                                           .arlock
		.UABChip_0_axi4_mmio_master_arcache               (uabchip_0_axi4_mmio_master_arcache),            //                                           .arcache
		.UABChip_0_axi4_mmio_master_arprot                (uabchip_0_axi4_mmio_master_arprot),             //                                           .arprot
		.UABChip_0_axi4_mmio_master_arqos                 (uabchip_0_axi4_mmio_master_arqos),              //                                           .arqos
		.UABChip_0_axi4_mmio_master_arvalid               (uabchip_0_axi4_mmio_master_arvalid),            //                                           .arvalid
		.UABChip_0_axi4_mmio_master_arready               (uabchip_0_axi4_mmio_master_arready),            //                                           .arready
		.UABChip_0_axi4_mmio_master_rid                   (uabchip_0_axi4_mmio_master_rid),                //                                           .rid
		.UABChip_0_axi4_mmio_master_rdata                 (uabchip_0_axi4_mmio_master_rdata),              //                                           .rdata
		.UABChip_0_axi4_mmio_master_rresp                 (uabchip_0_axi4_mmio_master_rresp),              //                                           .rresp
		.UABChip_0_axi4_mmio_master_rlast                 (uabchip_0_axi4_mmio_master_rlast),              //                                           .rlast
		.UABChip_0_axi4_mmio_master_rvalid                (uabchip_0_axi4_mmio_master_rvalid),             //                                           .rvalid
		.UABChip_0_axi4_mmio_master_rready                (uabchip_0_axi4_mmio_master_rready),             //                                           .rready
		.clk_clk_clk                                      (clk_clk),                                       //                                    clk_clk.clk
		.onchip_memory_reset1_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // onchip_memory_reset1_reset_bridge_in_reset.reset
		.UABChip_0_reset_reset_bridge_in_reset_reset      (uabchip_reset_reset),                           //      UABChip_0_reset_reset_bridge_in_reset.reset
		.onchip_memory_s1_address                         (mm_interconnect_1_onchip_memory_s1_address),    //                           onchip_memory_s1.address
		.onchip_memory_s1_write                           (mm_interconnect_1_onchip_memory_s1_write),      //                                           .write
		.onchip_memory_s1_readdata                        (mm_interconnect_1_onchip_memory_s1_readdata),   //                                           .readdata
		.onchip_memory_s1_writedata                       (mm_interconnect_1_onchip_memory_s1_writedata),  //                                           .writedata
		.onchip_memory_s1_byteenable                      (mm_interconnect_1_onchip_memory_s1_byteenable), //                                           .byteenable
		.onchip_memory_s1_chipselect                      (mm_interconnect_1_onchip_memory_s1_chipselect), //                                           .chipselect
		.onchip_memory_s1_clken                           (mm_interconnect_1_onchip_memory_s1_clken),      //                                           .clken
		.pio_0_s1_address                                 (mm_interconnect_1_pio_0_s1_address),            //                                   pio_0_s1.address
		.pio_0_s1_write                                   (mm_interconnect_1_pio_0_s1_write),              //                                           .write
		.pio_0_s1_readdata                                (mm_interconnect_1_pio_0_s1_readdata),           //                                           .readdata
		.pio_0_s1_writedata                               (mm_interconnect_1_pio_0_s1_writedata),          //                                           .writedata
		.pio_0_s1_chipselect                              (mm_interconnect_1_pio_0_s1_chipselect)          //                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~ddr3_h2f_reset_reset),              // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~ddr3_h2f_reset_reset),              // reset_in0.reset
		.clk            (mem_pll_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
